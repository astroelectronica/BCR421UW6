.title KiCad schematic
.include "C:/AE/BCR421UW6/BCR421UW6.spice.txt"
.include "C:/AE/BCR421UW6/SML-011VT_SPICE.lib"
D3 /LD2 /LD3 SML-011VT
D4 /LD3 /LD4 SML-011VT
R1 0 /REXT {REXT}
D1 VCC /LD1 SML-011VT
D2 /LD1 /LD2 SML-011VT
XU1 /EN /LD4 /LD4 0 /LD4 /REXT BCR421UW6
V2 /EN 0 DC PULSE(0 {VPUL} {DELAY} {TR} {TF} {DUTY} {CYCLE} 
V1 VCC 0 DC {VSOURCE} 
.end
