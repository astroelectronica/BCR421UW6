.title KiCad schematic
.include "C:/AE/BCR421UW6/BCR421UW6.spice.txt"
.include "C:/AE/BCR421UW6/SML-011VT_SPICE.lib"
D2 /LD1 /LD2 SML-011VT
D1 VCC /LD1 SML-011VT
V2 /EN 0 DC {EN} 
V1 VCC 0 DC {VSOURCE} 
D3 /LD2 /LD3 SML-011VT
D4 /LD3 /LD4 SML-011VT
R1 0 /REXT {REXT}
XU1 /EN /LD4 /LD4 0 /LD4 /REXT BCR421UW6
.end
